`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2018 10:21:50 PM
// Design Name: 
// Module Name: mux2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2_2
    #(parameter WIDTH = 32)
    (input logic [WIDTH-1:0] d0, d1,
     input logic [1:0] s,
     output logic [WIDTH-1:0] y);

assign y = ((s==2'b01)||(s==2'b10)||(s==2'b11) )? d1 : d0;

endmodule
