`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/07/2018 10:10:33 PM
// Design Name: 
// Module Name: Controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Controller(
    
    //Input
    input logic [6:0] Opcode, //7-bit opcode field from the instruction
    
    //Outputs
    output logic ALUSrc,//0: The second ALU operand comes from the second register file output (Read data 2); 
                  //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic MemtoReg, //0: The value fed to the register Write data input comes from the ALU.
                     //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input 
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic Branch,  //0: branch is not taken; 1: branch is taken
    output logic [1:0] ALUOp,
    output logic [1:0] PC_Reg
);

//    localparam R_TYPE = 7'b0110011;
//    localparam LW     = 7'b0000011;
//    localparam SW     = 7'b0100011;
//    localparam BR     = 7'b1100011;
//    localparam RTypeI = 7'b0010011; //addi,ori,andi
    
    logic [6:0] LUI,AUIPC,JAL,JALR,B_TYPE,R_TYPE, LW, SW, RTypeI;
    

    assign  LUI    = 7'b0110111;
    assign  AUIPC  = 7'b0010111;

    assign  JAL    = 7'b1101111;
    assign  JALR   = 7'b1100111;

    assign  B_TYPE = 7'b1100011;

    assign  R_TYPE = 7'b0110011;
    assign  LW     = 7'b0000011;
    assign  SW     = 7'b0100011;
    assign  RTypeI = 7'b0010011; //addi,ori,andi

// ALUOp indicates whether the operation to be performed should be add (00) for loads and stores, 
// subtract and test if zero (01) for beq,
// or be determined by the operation encoded in the funct7 and funct3 fields (10).


  assign ALUSrc   = (Opcode==LW || Opcode==SW || Opcode == RTypeI || Opcode == LUI );
  assign MemtoReg = (Opcode==LW);
  assign RegWrite = (Opcode==R_TYPE || Opcode==LW || Opcode == RTypeI || Opcode == LUI || Opcode == AUIPC || Opcode == JALR || Opcode ==JAL );
  assign MemRead  = (Opcode==LW);
  assign MemWrite = (Opcode==SW);
  assign Branch = (Opcode==B_TYPE || Opcode == JAL );
  
  //Need to be modified 
  assign ALUOp =  Opcode == B_TYPE ? 2'b01:(Opcode == R_TYPE? 2'b10:(Opcode == RTypeI ? 2'b11:2'b00));
  //Additional Mux added
  assign PC_Reg = Opcode == AUIPC? 2'b01:(Opcode == JAL? 2'b10:(Opcode == JALR ? 2'b11:2'b00));
  

endmodule
